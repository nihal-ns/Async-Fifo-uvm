`define ASIZE 8
`define DSIZE 4
